-- Cosine table signal
-- 1250 values in table represents as 11 bit bin number "angle"
-- Each values is 7 bit number from 111001 (77) to 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity cos_table_gen is
    port (
        clk : in std_logic;
        reset : in std_logic;
        cosine_out : out std_logic_vector(6 downto 0)
    );
end entity cos_table_gen;

architecture src of cos_table_gen is

    signal angle : std_logic_vector(10 downto 0) := (others => '0');
  
    type cosine_table_type is array (0 to 1249) of std_logic_vector(6 downto 0);
    
    constant cosine_table : cosine_table_type := (
        "1111001", -- 77
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111001",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1111000",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110111",
        "1110110",
        "1110110",
        "1110110",
        "1110110",
        "1110110",
        "1110110",
        "1110110",
        "1110110",
        "1110110",
        "1110110",
        "1110110",
        "1110110",
        "1110110",
        "1110110",
        "1110110",
        "1110110",
        "1110110",
        "1110110",
        "1110110",
        "1110110",
        "1110110",
        "1110101",
        "1110101",
        "1110101",
        "1110101",
        "1110101",
        "1110101",
        "1110101",
        "1110101",
        "1110101",
        "1110101",
        "1110101",
        "1110101",
        "1110101",
        "1110101",
        "1110101",
        "1110101",
        "1110101",
        "1110101",
        "1110101",
        "1110100",
        "1110100",
        "1110100",
        "1110100",
        "1110100",
        "1110100",
        "1110100",
        "1110100",
        "1110100",
        "1110100",
        "1110100",
        "1110100",
        "1110100",
        "1110100",
        "1110100",
        "1110100",
        "1110011",
        "1110011",
        "1110011",
        "1110011",
        "1110011",
        "1110011",
        "1110011",
        "1110011",
        "1110011",
        "1110011",
        "1110011",
        "1110011",
        "1110011",
        "1110011",
        "1110011",
        "1110011",
        "1110010",
        "1110010",
        "1110010",
        "1110010",
        "1110010",
        "1110010",
        "1110010",
        "1110010",
        "1110010",
        "1110010",
        "1110010",
        "1110010",
        "1110010",
        "1110010",
        "1110001",
        "1110001",
        "1110001",
        "1110001",
        "1110001",
        "1110001",
        "1110001",
        "1110001",
        "1110001",
        "1110001",
        "1110001",
        "1110001",
        "1110001",
        "1110001",
        "1110000",
        "1110000",
        "1110000",
        "1110000",
        "1110000",
        "1110000",
        "1110000",
        "1110000",
        "1110000",
        "1110000",
        "1110000",
        "1110000",
        "1110000",
        "1101111",
        "1101111",
        "1101111",
        "1101111",
        "1101111",
        "1101111",
        "1101111",
        "1101111",
        "1101111",
        "1101111",
        "1101111",
        "1101111",
        "1101110",
        "1101110",
        "1101110",
        "1101110",
        "1101110",
        "1101110",
        "1101110",
        "1101110",
        "1101110",
        "1101110",
        "1101110",
        "1101101",
        "1101101",
        "1101101",
        "1101101",
        "1101101",
        "1101101",
        "1101101",
        "1101101",
        "1101101",
        "1101101",
        "1101101",
        "1101101",
        "1101100",
        "1101100",
        "1101100",
        "1101100",
        "1101100",
        "1101100",
        "1101100",
        "1101100",
        "1101100",
        "1101100",
        "1101100",
        "1101011",
        "1101011",
        "1101011",
        "1101011",
        "1101011",
        "1101011",
        "1101011",
        "1101011",
        "1101011",
        "1101011",
        "1101010",
        "1101010",
        "1101010",
        "1101010",
        "1101010",
        "1101010",
        "1101010",
        "1101010",
        "1101010",
        "1101010",
        "1101001",
        "1101001",
        "1101001",
        "1101001",
        "1101001",
        "1101001",
        "1101001",
        "1101001",
        "1101001",
        "1101001",
        "1101000",
        "1101000",
        "1101000",
        "1101000",
        "1101000",
        "1101000",
        "1101000",
        "1101000",
        "1101000",
        "1101000",
        "1100111",
        "1100111",
        "1100111",
        "1100111",
        "1100111",
        "1100111",
        "1100111",
        "1100111",
        "1100111",
        "1100111",
        "1100110",
        "1100110",
        "1100110",
        "1100110",
        "1100110",
        "1100110",
        "1100110",
        "1100110",
        "1100110",
        "1100101",
        "1100101",
        "1100101",
        "1100101",
        "1100101",
        "1100101",
        "1100101",
        "1100101",
        "1100101",
        "1100100",
        "1100100",
        "1100100",
        "1100100",
        "1100100",
        "1100100",
        "1100100",
        "1100100",
        "1100100",
        "1100011",
        "1100011",
        "1100011",
        "1100011",
        "1100011",
        "1100011",
        "1100011",
        "1100011",
        "1100011",
        "1100010",
        "1100010",
        "1100010",
        "1100010",
        "1100010",
        "1100010",
        "1100010",
        "1100010",
        "1100001",
        "1100001",
        "1100001",
        "1100001",
        "1100001",
        "1100001",
        "1100001",
        "1100001",
        "1100001",
        "1100000",
        "1100000",
        "1100000",
        "1100000",
        "1100000",
        "1100000",
        "1100000",
        "1100000",
        "1011111",
        "1011111",
        "1011111",
        "1011111",
        "1011111",
        "1011111",
        "1011111",
        "1011111",
        "1011110",
        "1011110",
        "1011110",
        "1011110",
        "1011110",
        "1011110",
        "1011110",
        "1011110",
        "1011110",
        "1011101",
        "1011101",
        "1011101",
        "1011101",
        "1011101",
        "1011101",
        "1011101",
        "1011101",
        "1011100",
        "1011100",
        "1011100",
        "1011100",
        "1011100",
        "1011100",
        "1011100",
        "1011100",
        "1011011",
        "1011011",
        "1011011",
        "1011011",
        "1011011",
        "1011011",
        "1011011",
        "1011010",
        "1011010",
        "1011010",
        "1011010",
        "1011010",
        "1011010",
        "1011010",
        "1011010",
        "1011001",
        "1011001",
        "1011001",
        "1011001",
        "1011001",
        "1011001",
        "1011001",
        "1011001",
        "1011000",
        "1011000",
        "1011000",
        "1011000",
        "1011000",
        "1011000",
        "1011000",
        "1011000",
        "1010111",
        "1010111",
        "1010111",
        "1010111",
        "1010111",
        "1010111",
        "1010111",
        "1010110",
        "1010110",
        "1010110",
        "1010110",
        "1010110",
        "1010110",
        "1010110",
        "1010110",
        "1010101",
        "1010101",
        "1010101",
        "1010101",
        "1010101",
        "1010101",
        "1010101",
        "1010100",
        "1010100",
        "1010100",
        "1010100",
        "1010100",
        "1010100",
        "1010100",
        "1010011",
        "1010011",
        "1010011",
        "1010011",
        "1010011",
        "1010011",
        "1010011",
        "1010011",
        "1010010",
        "1010010",
        "1010010",
        "1010010",
        "1010010",
        "1010010",
        "1010010",
        "1010001",
        "1010001",
        "1010001",
        "1010001",
        "1010001",
        "1010001",
        "1010001",
        "1010000",
        "1010000",
        "1010000",
        "1010000",
        "1010000",
        "1010000",
        "1010000",
        "1010000",
        "1001111",
        "1001111",
        "1001111",
        "1001111",
        "1001111",
        "1001111",
        "1001111",
        "1001110",
        "1001110",
        "1001110",
        "1001110",
        "1001110",
        "1001110",
        "1001110",
        "1001101",
        "1001101",
        "1001101",
        "1001101",
        "1001101",
        "1001101",
        "1001101",
        "1001100",
        "1001100",
        "1001100",
        "1001100",
        "1001100",
        "1001100",
        "1001100",
        "1001011",
        "1001011",
        "1001011",
        "1001011",
        "1001011",
        "1001011",
        "1001011",
        "1001010",
        "1001010",
        "1001010",
        "1001010",
        "1001010",
        "1001010",
        "1001010",
        "1001001",
        "1001001",
        "1001001",
        "1001001",
        "1001001",
        "1001001",
        "1001001",
        "1001000",
        "1001000",
        "1001000",
        "1001000",
        "1001000",
        "1001000",
        "1001000",
        "1000111",
        "1000111",
        "1000111",
        "1000111",
        "1000111",
        "1000111",
        "1000111",
        "1000110",
        "1000110",
        "1000110",
        "1000110",
        "1000110",
        "1000110",
        "1000110",
        "1000101",
        "1000101",
        "1000101",
        "1000101",
        "1000101",
        "1000101",
        "1000101",
        "1000100",
        "1000100",
        "1000100",
        "1000100",
        "1000100",
        "1000100",
        "1000100",
        "1000011",
        "1000011",
        "1000011",
        "1000011",
        "1000011",
        "1000011",
        "1000011",
        "1000010",
        "1000010",
        "1000010",
        "1000010",
        "1000010",
        "1000010",
        "1000010",
        "1000001",
        "1000001",
        "1000001",
        "1000001",
        "1000001",
        "1000001",
        "1000001",
        "1000000",
        "1000000",
        "1000000",
        "1000000",
        "1000000",
        "1000000",
        "1000000",
        "0111111",
        "0111111",
        "0111111",
        "0111111",
        "0111111",
        "0111111",
        "0111110",
        "0111110",
        "0111110",
        "0111110",
        "0111110",
        "0111110",
        "0111110",
        "0111101",
        "0111101",
        "0111101",
        "0111101",
        "0111101",
        "0111101",
        "0111101",
        "0111100",
        "0111100",
        "0111100",
        "0111100",
        "0111100",
        "0111100",
        "0111100",
        "0111011",
        "0111011",
        "0111011",
        "0111011",
        "0111011",
        "0111011",
        "0111011",
        "0111010",
        "0111010",
        "0111010",
        "0111010",
        "0111010",
        "0111010",
        "0111010",
        "0111001",
        "0111001",
        "0111001",
        "0111001",
        "0111001",
        "0111001",
        "0111001",
        "0111000",
        "0111000",
        "0111000",
        "0111000",
        "0111000",
        "0111000",
        "0111000",
        "0110111",
        "0110111",
        "0110111",
        "0110111",
        "0110111",
        "0110111",
        "0110111",
        "0110110",
        "0110110",
        "0110110",
        "0110110",
        "0110110",
        "0110110",
        "0110110",
        "0110101",
        "0110101",
        "0110101",
        "0110101",
        "0110101",
        "0110101",
        "0110101",
        "0110100",
        "0110100",
        "0110100",
        "0110100",
        "0110100",
        "0110100",
        "0110100",
        "0110011",
        "0110011",
        "0110011",
        "0110011",
        "0110011",
        "0110011",
        "0110011",
        "0110010",
        "0110010",
        "0110010",
        "0110010",
        "0110010",
        "0110010",
        "0110010",
        "0110001",
        "0110001",
        "0110001",
        "0110001",
        "0110001",
        "0110001",
        "0110001",
        "0110000",
        "0110000",
        "0110000",
        "0110000",
        "0110000",
        "0110000",
        "0110000",
        "0110000",
        "0101111",
        "0101111",
        "0101111",
        "0101111",
        "0101111",
        "0101111",
        "0101111",
        "0101110",
        "0101110",
        "0101110",
        "0101110",
        "0101110",
        "0101110",
        "0101110",
        "0101101",
        "0101101",
        "0101101",
        "0101101",
        "0101101",
        "0101101",
        "0101101",
        "0101100",
        "0101100",
        "0101100",
        "0101100",
        "0101100",
        "0101100",
        "0101100",
        "0101100",
        "0101011",
        "0101011",
        "0101011",
        "0101011",
        "0101011",
        "0101011",
        "0101011",
        "0101010",
        "0101010",
        "0101010",
        "0101010",
        "0101010",
        "0101010",
        "0101010",
        "0101001",
        "0101001",
        "0101001",
        "0101001",
        "0101001",
        "0101001",
        "0101001",
        "0101001",
        "0101000",
        "0101000",
        "0101000",
        "0101000",
        "0101000",
        "0101000",
        "0101000",
        "0101000",
        "0100111",
        "0100111",
        "0100111",
        "0100111",
        "0100111",
        "0100111",
        "0100111",
        "0100110",
        "0100110",
        "0100110",
        "0100110",
        "0100110",
        "0100110",
        "0100110",
        "0100110",
        "0100101",
        "0100101",
        "0100101",
        "0100101",
        "0100101",
        "0100101",
        "0100101",
        "0100101",
        "0100100",
        "0100100",
        "0100100",
        "0100100",
        "0100100",
        "0100100",
        "0100100",
        "0100011",
        "0100011",
        "0100011",
        "0100011",
        "0100011",
        "0100011",
        "0100011",
        "0100011",
        "0100010",
        "0100010",
        "0100010",
        "0100010",
        "0100010",
        "0100010",
        "0100010",
        "0100010",
        "0100001",
        "0100001",
        "0100001",
        "0100001",
        "0100001",
        "0100001",
        "0100001",
        "0100001",
        "0100001",
        "0100000",
        "0100000",
        "0100000",
        "0100000",
        "0100000",
        "0100000",
        "0100000",
        "0100000",
        "0011111",
        "0011111",
        "0011111",
        "0011111",
        "0011111",
        "0011111",
        "0011111",
        "0011111",
        "0011110",
        "0011110",
        "0011110",
        "0011110",
        "0011110",
        "0011110",
        "0011110",
        "0011110",
        "0011110",
        "0011101",
        "0011101",
        "0011101",
        "0011101",
        "0011101",
        "0011101",
        "0011101",
        "0011101",
        "0011100",
        "0011100",
        "0011100",
        "0011100",
        "0011100",
        "0011100",
        "0011100",
        "0011100",
        "0011100",
        "0011011",
        "0011011",
        "0011011",
        "0011011",
        "0011011",
        "0011011",
        "0011011",
        "0011011",
        "0011011",
        "0011010",
        "0011010",
        "0011010",
        "0011010",
        "0011010",
        "0011010",
        "0011010",
        "0011010",
        "0011010",
        "0011001",
        "0011001",
        "0011001",
        "0011001",
        "0011001",
        "0011001",
        "0011001",
        "0011001",
        "0011001",
        "0011000",
        "0011000",
        "0011000",
        "0011000",
        "0011000",
        "0011000",
        "0011000",
        "0011000",
        "0011000",
        "0011000",
        "0010111",
        "0010111",
        "0010111",
        "0010111",
        "0010111",
        "0010111",
        "0010111",
        "0010111",
        "0010111",
        "0010111",
        "0010110",
        "0010110",
        "0010110",
        "0010110",
        "0010110",
        "0010110",
        "0010110",
        "0010110",
        "0010110",
        "0010110",
        "0010101",
        "0010101",
        "0010101",
        "0010101",
        "0010101",
        "0010101",
        "0010101",
        "0010101",
        "0010101",
        "0010101",
        "0010100",
        "0010100",
        "0010100",
        "0010100",
        "0010100",
        "0010100",
        "0010100",
        "0010100",
        "0010100",
        "0010100",
        "0010011",
        "0010011",
        "0010011",
        "0010011",
        "0010011",
        "0010011",
        "0010011",
        "0010011",
        "0010011",
        "0010011",
        "0010011",
        "0010010",
        "0010010",
        "0010010",
        "0010010",
        "0010010",
        "0010010",
        "0010010",
        "0010010",
        "0010010",
        "0010010",
        "0010010",
        "0010010",
        "0010001",
        "0010001",
        "0010001",
        "0010001",
        "0010001",
        "0010001",
        "0010001",
        "0010001",
        "0010001",
        "0010001",
        "0010001",
        "0010000",
        "0010000",
        "0010000",
        "0010000",
        "0010000",
        "0010000",
        "0010000",
        "0010000",
        "0010000",
        "0010000",
        "0010000",
        "0010000",
        "0001111",
        "0001111",
        "0001111",
        "0001111",
        "0001111",
        "0001111",
        "0001111",
        "0001111",
        "0001111",
        "0001111",
        "0001111",
        "0001111",
        "0001111",
        "0001110",
        "0001110",
        "0001110",
        "0001110",
        "0001110",
        "0001110",
        "0001110",
        "0001110",
        "0001110",
        "0001110",
        "0001110",
        "0001110",
        "0001110",
        "0001110",
        "0001101",
        "0001101",
        "0001101",
        "0001101",
        "0001101",
        "0001101",
        "0001101",
        "0001101",
        "0001101",
        "0001101",
        "0001101",
        "0001101",
        "0001101",
        "0001101",
        "0001100",
        "0001100",
        "0001100",
        "0001100",
        "0001100",
        "0001100",
        "0001100",
        "0001100",
        "0001100",
        "0001100",
        "0001100",
        "0001100",
        "0001100",
        "0001100",
        "0001100",
        "0001100",
        "0001011",
        "0001011",
        "0001011",
        "0001011",
        "0001011",
        "0001011",
        "0001011",
        "0001011",
        "0001011",
        "0001011",
        "0001011",
        "0001011",
        "0001011",
        "0001011",
        "0001011",
        "0001011",
        "0001010",
        "0001010",
        "0001010",
        "0001010",
        "0001010",
        "0001010",
        "0001010",
        "0001010",
        "0001010",
        "0001010",
        "0001010",
        "0001010",
        "0001010",
        "0001010",
        "0001010",
        "0001010",
        "0001010",
        "0001010",
        "0001010",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001001",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0001000",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000111",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110",
        "0000110"
    );

    signal angle_reg : std_logic_vector(10 downto 0);
    signal cosine_value : std_logic_vector(6 downto 0);
    
begin
    read_table : process(clk, reset, angle)
    begin
        if reset = '1' then
            angle_reg <= (others => '0');
            cosine_value <= (others => '0');
        elsif rising_edge(clk) then
            angle_reg <= angle;
            cosine_value <= cosine_table(to_integer(unsigned(angle_reg)));
        end if;
    end process;
    
    cosine_out <= cosine_value;
    
    angle_generator : process(clk, angle)
        variable angle_reset : std_logic := '0';
        variable angle_updown : std_logic := '0';
    begin
        if rising_edge(clk) then
            if angle_reset = '1' then
                angle <= b"00000000000";
                angle_updown := '1';
            elsif angle_updown = '1' and angle < b"10011100001" then
                angle <= std_logic_vector(unsigned(angle) + b"00000000001");
            elsif angle_updown = '0' and angle > b"00000000000" then
                angle <= std_logic_vector(unsigned(angle) - b"00000000001");
            elsif angle = b"00000000000" then
                angle_updown := '1';
                angle <= std_logic_vector(unsigned(angle) + b"00000000001");
            elsif angle = b"10011100001" then
                angle_updown := '0';
                angle <= std_logic_vector(unsigned(angle) - b"00000000001");
            end if;
        end if;
    end process;

end src;